library verilog;
use verilog.vl_types.all;
entity lab3_p1_vlg_vec_tst is
end lab3_p1_vlg_vec_tst;
