library verilog;
use verilog.vl_types.all;
entity Lab3_p2_vlg_check_tst is
    port(
        f0              : in     vl_logic;
        f1              : in     vl_logic;
        f2              : in     vl_logic;
        f3              : in     vl_logic;
        f4              : in     vl_logic;
        f5              : in     vl_logic;
        f6              : in     vl_logic;
        f7              : in     vl_logic;
        f8              : in     vl_logic;
        f9              : in     vl_logic;
        f10             : in     vl_logic;
        f11             : in     vl_logic;
        f12             : in     vl_logic;
        f13             : in     vl_logic;
        f14             : in     vl_logic;
        f15             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab3_p2_vlg_check_tst;
