library verilog;
use verilog.vl_types.all;
entity lab3_p1_vlg_check_tst is
    port(
        F0              : in     vl_logic;
        F1              : in     vl_logic;
        F2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab3_p1_vlg_check_tst;
