library verilog;
use verilog.vl_types.all;
entity Lab3_p2 is
    port(
        f15             : out    vl_logic;
        W               : in     vl_logic;
        X               : in     vl_logic;
        Y               : in     vl_logic;
        Z               : in     vl_logic;
        f14             : out    vl_logic;
        f13             : out    vl_logic;
        f12             : out    vl_logic;
        f11             : out    vl_logic;
        f10             : out    vl_logic;
        f9              : out    vl_logic;
        f8              : out    vl_logic;
        f7              : out    vl_logic;
        f6              : out    vl_logic;
        f5              : out    vl_logic;
        f4              : out    vl_logic;
        f3              : out    vl_logic;
        f2              : out    vl_logic;
        f1              : out    vl_logic;
        f0              : out    vl_logic
    );
end Lab3_p2;
