library verilog;
use verilog.vl_types.all;
entity lab6_p2 is
    port(
        A               : out    vl_logic;
        A2              : in     vl_logic;
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        A3              : in     vl_logic;
        b               : out    vl_logic;
        c               : out    vl_logic;
        d               : out    vl_logic;
        e               : out    vl_logic;
        f               : out    vl_logic;
        g               : out    vl_logic
    );
end lab6_p2;
