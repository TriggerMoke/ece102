library verilog;
use verilog.vl_types.all;
entity lab3_p1 is
    port(
        F2              : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        F1              : out    vl_logic;
        F0              : out    vl_logic
    );
end lab3_p1;
